

module base_project (
  output LED0,
  input test_pin
);

assign LED0 = test_pin;

endmodule
